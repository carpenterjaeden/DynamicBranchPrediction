module XOR ( input a, input b, output out);
    assign out = a ^ b; // ^ is the XOR operator
endmodule