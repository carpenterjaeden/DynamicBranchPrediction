module Branch_Predictor(
);

endmodule